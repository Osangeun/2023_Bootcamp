library verilog;
use verilog.vl_types.all;
entity tb_johnson_cnt is
end tb_johnson_cnt;
