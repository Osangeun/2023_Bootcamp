library verilog;
use verilog.vl_types.all;
entity tb_D_FF is
end tb_D_FF;
