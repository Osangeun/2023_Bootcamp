library verilog;
use verilog.vl_types.all;
entity tb_binary_cnt is
end tb_binary_cnt;
