library verilog;
use verilog.vl_types.all;
entity tb_ring_cnt is
end tb_ring_cnt;
