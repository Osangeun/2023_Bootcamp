library verilog;
use verilog.vl_types.all;
entity ring_cnt is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        q               : out    vl_logic_vector(3 downto 0)
    );
end ring_cnt;
